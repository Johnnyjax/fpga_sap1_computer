library verilog;
use verilog.vl_types.all;
entity sap_1_vlg_vec_tst is
end sap_1_vlg_vec_tst;
